LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY Controller IS
	PORT (
		opcode : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		reset_input : IN STD_LOGIC;
		ZF : IN STD_LOGIC;
		jump, jumpZ, rst, immEnable, immFlush, memoryWrite, memoryRead, returnEnable, callEnable, aluImm, writeEnable, alu_enable, oneoperand, swap_enable, protect_enable, free_enable, push_enable, pop_enable, Out_port : OUT STD_LOGIC;
		opcode_to_alu : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		INT, RTI : OUT STD_LOGIC
	);
END Controller;

ARCHITECTURE controller_model OF Controller IS
BEGIN
	PROCESS (opcode, reset_input)
	BEGIN
		IF reset_input = '1' THEN
			rst <= '1';
			jump <= '0';
			jumpZ <= '0';
			immEnable <= '0';
			immFlush <= '0';
			memoryWrite <= '0';
			memoryRead <= '0';
			returnEnable <= '0';
			callEnable <= '0';
			aluImm <= '0';
			writeEnable <= '0';
			alu_enable <= '0';
			oneoperand <= '0';
			INT <= '0';
			RTI <= '0';
			protect_enable <= '0';
			free_enable <= '0';
			push_enable <= '0';
			pop_enable <= '0';
			Out_port <= '0';
		ELSE
			CASE opcode IS
				WHEN "0000000" =>
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '0';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '0';
					alu_enable <= '0';
					oneoperand <= '0';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "0000001" => --reset
					rst <= '1';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '0';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '0';
					alu_enable <= '0';
					oneoperand <= '0';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "0101001" => -- SWAP
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '0';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '1';
					swap_enable <= '1';
					alu_enable <= '0';
					oneoperand <= '0';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "0101000" => --move
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '0';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '1';
					swap_enable <= '0';
					alu_enable <= '0';
					oneoperand <= '0';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "0001101" => --in
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '0';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '1';
					alu_enable <= '0';
					oneoperand <= '1';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "0110000" | "0110001" | "0110010" | "0110011" | "0110100" => --add|sub|and|or|xor
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '0';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '1';
					alu_enable <= '1';
					oneoperand <= '0';
					INT <= '0';
					RTI <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					protect_enable <= '0';
					Out_port <= '0';
				WHEN "0001011" | "0001010" | "0001001" | "0001000" => --dec|inc|neg|not
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '0';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '1';
					alu_enable <= '1';
					oneoperand <= '1';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "0001100" => --out
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '0';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '0';
					alu_enable <= '0';
					oneoperand <= '0';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '1';
				WHEN "0100000" => --cmp
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '0';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '0';
					alu_enable <= '1';
					oneoperand <= '0';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "0111000" | "0111001" => --addi|subi
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '1';
					immFlush <= '1';
					memoryWrite <= '0';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '1';
					writeEnable <= '1';
					alu_enable <= '1';
					oneoperand <= '0';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "1001000" => --push
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '1';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '0';
					alu_enable <= '0';
					oneoperand <= '1';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '1';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "1001001" => --pop
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '0';
					memoryRead <= '1';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '1';
					alu_enable <= '0';
					oneoperand <= '1';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '1';
					Out_port <= '0';
				WHEN "1010000" => --Load immediate
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '1';
					immFlush <= '1';
					memoryWrite <= '0';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '1';
					writeEnable <= '1';
					alu_enable <= '0';
					oneoperand <= '0';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "1011000" => --Load
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '1';
					immFlush <= '1';
					memoryWrite <= '0';
					memoryRead <= '1';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '1';
					alu_enable <= '0';
					oneoperand <= '0';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "1011001" => --store
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '1';
					immFlush <= '1';
					memoryWrite <= '1';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '1';
					writeEnable <= '0';
					alu_enable <= '1';
					oneoperand <= '0';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "1101000" => --jz
					rst <= '0';
					jump <= '0';
					jumpZ <= ZF;
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '0';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '0';
					alu_enable <= '1';
					oneoperand <= '1';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "1101001" => --jump
					rst <= '0';
					jump <= '1';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '0';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '0';
					alu_enable <= '0';
					oneoperand <= '1';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "1101010" => --call
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '1';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '1';
					aluImm <= '0';
					writeEnable <= '0';
					alu_enable <= '0';
					oneoperand <= '1';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "1100000" => --return
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '0';
					memoryRead <= '1';
					returnEnable <= '1';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '0';
					alu_enable <= '0';
					oneoperand <= '0';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "0000010" => -- INT
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '1';
					memoryRead <= '1';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '0';
					alu_enable <= '0';
					oneoperand <= '0';
					INT <= '1';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "1100001" => -- RTI
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '0';
					memoryRead <= '1';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '0';
					alu_enable <= '0';
					oneoperand <= '0';
					INT <= '0';
					RTI <= '1';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "1000000" => -- PROTECT
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '1';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '0';
					alu_enable <= '0';
					oneoperand <= '0';
					INT <= '0';
					RTI <= '1';
					protect_enable <= '1';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN "1000001" => -- FREE
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '1';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '0';
					alu_enable <= '0';
					oneoperand <= '0';
					INT <= '0';
					RTI <= '1';
					protect_enable <= '1';
					free_enable <= '1';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
				WHEN OTHERS =>
					rst <= '0';
					jump <= '0';
					jumpZ <= '0';
					immEnable <= '0';
					immFlush <= '0';
					memoryWrite <= '0';
					memoryRead <= '0';
					returnEnable <= '0';
					callEnable <= '0';
					aluImm <= '0';
					writeEnable <= '0';
					alu_enable <= '0';
					oneoperand <= '0';
					INT <= '0';
					RTI <= '0';
					protect_enable <= '0';
					free_enable <= '0';
					push_enable <= '0';
					pop_enable <= '0';
					Out_port <= '0';
			END CASE;
		END IF;
		opcode_to_alu <= opcode;
	END PROCESS;
END ARCHITECTURE;