LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY CCR IS
    PORT (
        CCR_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        CCR_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END CCR;

ARCHITECTURE BEHAVIOR OF CCR IS
BEGIN
    CCR_OUT <= CCR_IN;
END ARCHITECTURE;